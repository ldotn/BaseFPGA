`timescale 1 ps / 1 ps

module cache_testbed;
	
	Read_Only_Cache cache;
	
endmodule