`timescale 1 ps / 1 ps

module Cache_Testbench;
	
	Read_Only_Cache cache;
	
endmodule